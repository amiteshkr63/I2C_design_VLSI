`define DATA_WIDTH 8
`define ADDR_WIDTH 7